`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/26/2024 05:36:00 PM
// Design Name: 
// Module Name: top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module top(
	input              APB_hbm_reset,
	input              HBM_REF_CLK_0,
    input             APB_0_PCLK,
    input             AXI_ACLK,                                  // Clock signal
    input             AXI_ARESET_N,                                  // Reset signal
	input write_enable [16],
	input read_enable [16],
	input [255:0] write_data [16],
	input [33:0] write_address [16],
	input [33:0] read_address [16]	

    );

    logic [33:0] AXI_ARADDR [16];            // Read data addresses
    logic [1:0] AXI_ARBURST [16];            // Read burst types
    logic [5:0] AXI_ARID [16];               // Read IDs
    logic [3:0] AXI_ARLEN [16];              // Read transfer lengths
    logic [2:0] AXI_ARSIZE [16];             // Read transfer sizes
    logic AXI_ARVALID [16];                  // Read address valid signals
    logic [33:0] AXI_AWADDR [16];            // Write data addresses
    logic [1:0] AXI_AWBURST [16];            // Write burst types
    logic [5:0] AXI_AWID [16];               // Write IDs
    logic [3:0] AXI_AWLEN [16];              // Write transfer lengths
    logic [2:0] AXI_AWSIZE [16];             // Write transfer sizes
    logic AXI_AWVALID [16];                  // Write address valid signals
    logic AXI_RREADY [16];                   // Read response ready signals
    logic AXI_BREADY [16];                   // Write response ready signals
    logic [255:0] AXI_WDATA [16];             // Write data
    logic [31:0] AXI_WSTRB [16];              // Write byte enables
    logic AXI_WLAST [16];                    // Write last transfer cycles
    logic [31:0] AXI_WDATA_PARITY [16];             // Write data parity
    logic  AXI_WVALID [16];                   // Write data valid signals	
    logic  AXI_ARREADY [16];                 // Read address ready signals
    logic  AXI_AWREADY [16];                 // Write address ready signals
	logic  AXI_WREADY [16];
    logic  [255:0] AXI_RDATA [16];            // Read data
    logic  [1:0] AXI_RRESP [16];             // Read responses
    logic  AXI_RLAST [16];                   // Read last transfer cycles
    logic  AXI_RVALID [16];                  // Read data valid signals
    logic  [5:0] AXI_RID [16];               // Read IDs
    logic  [5:0] AXI_BID [16];              // Write IDs
    logic  [1:0] AXI_BRESP [16];             // Write responses
    logic  AXI_BVALID [16];                   // Write data valid signals
	logic [31:0] AXI_RDATA_PARITY [16];             // Write data parity

	
axi_master_control_16 axi_master_control_16
(
    .AXI_ACLK(AXI_ACLK),
    .AXI_ARESET_N(AXI_ARESET_N),
    .AXI_ARADDR(AXI_ARADDR),
    .AXI_ARBURST(AXI_ARBURST),
    .AXI_ARID(AXI_ARID),
    .AXI_ARLEN(AXI_ARLEN),
    .AXI_ARSIZE(AXI_ARSIZE),
    .AXI_ARVALID(AXI_ARVALID),
    .AXI_AWADDR(AXI_AWADDR),
    .AXI_AWBURST(AXI_AWBURST),
    .AXI_AWID(AXI_AWID),
    .AXI_AWLEN(AXI_AWLEN),
    .AXI_AWSIZE(AXI_AWSIZE),
    .AXI_AWVALID(AXI_AWVALID),
    .AXI_RREADY(AXI_RREADY),
    .AXI_BREADY(AXI_BREADY),
    .AXI_WDATA(AXI_WDATA),
    .AXI_WSTRB(AXI_WSTRB),
    .AXI_WLAST(AXI_WLAST),
    .AXI_WDATA_PARITY(AXI_WDATA_PARITY),
    .AXI_WVALID(AXI_WVALID),
    .AXI_ARREADY(AXI_ARREADY),
    .AXI_AWREADY(AXI_AWREADY),
    .AXI_WREADY(AXI_WREADY),
    .AXI_RDATA(AXI_RDATA),
    .AXI_RRESP(AXI_RRESP),
    .AXI_RLAST(AXI_RLAST),
    .AXI_RVALID(AXI_RVALID),
    .AXI_RID(AXI_RID),
    .AXI_BID(AXI_BID),
    .AXI_BRESP(AXI_BRESP),
    .AXI_BVALID(AXI_BVALID),
    .write_enable(write_enable),
    .read_enable(read_enable),
    .write_data(write_data),
    .write_address(write_address),
    .read_address(read_address)
);

logic apb_complete_0;

logic    [ 31:0]  APB_0_PWDATA;
logic    [ 21:0]  APB_0_PADDR;
logic             APB_0_PENABLE;
logic             APB_0_PSEL;
logic             APB_0_PWRITE;
logic    [ 31:0]  APB_0_PRDATA;
logic             APB_0_PREADY;
logic             APB_0_PSLVERR;
always_comb APB_0_PADDR = '0;
always_comb APB_0_PENABLE = '0;
always_comb APB_0_PSEL = '0;
always_comb APB_0_PWDATA = '0;
always_comb APB_0_PWRITE = '0;

hbm_0 u_hbm_0
(
  .HBM_REF_CLK_0                 (HBM_REF_CLK_0)
  ,.AXI_00_ACLK                  (AXI_ACLK           )
  ,.AXI_00_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_00_ARADDR                (AXI_ARADDR[0]      )
  ,.AXI_00_ARBURST               (AXI_ARBURST[0]     )
  ,.AXI_00_ARID                  (AXI_ARID[0]        )
  ,.AXI_00_ARLEN                 (AXI_ARLEN[0]       )
  ,.AXI_00_ARSIZE                (AXI_ARSIZE[0]      )
  ,.AXI_00_ARVALID               (AXI_ARVALID[0]     )
  ,.AXI_00_AWADDR                (AXI_AWADDR[0]      )
  ,.AXI_00_AWBURST               (AXI_AWBURST[0]     )
  ,.AXI_00_AWID                  (AXI_AWID[0]        )
  ,.AXI_00_AWLEN                 (AXI_AWLEN[0]       )
  ,.AXI_00_AWSIZE                (AXI_AWSIZE[0]      )
  ,.AXI_00_AWVALID               (AXI_AWVALID[0]     )
  ,.AXI_00_RREADY                (AXI_RREADY[0]      )
  ,.AXI_00_BREADY                (AXI_BREADY[0]      )
  ,.AXI_00_WDATA                 (AXI_WDATA[0]       )
  ,.AXI_00_WLAST                 (AXI_WLAST[0]       )
  ,.AXI_00_WSTRB                 (AXI_WSTRB[0]       )
  ,.AXI_00_WDATA_PARITY          (AXI_WDATA_PARITY[0])
  ,.AXI_00_WVALID                (AXI_WVALID[0]      )
  ,.AXI_01_ACLK                  (AXI_ACLK           )
  ,.AXI_01_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_01_ARADDR                (AXI_ARADDR[1]      )
  ,.AXI_01_ARBURST               (AXI_ARBURST[1]     )
  ,.AXI_01_ARID                  (AXI_ARID[1]        )
  ,.AXI_01_ARLEN                 (AXI_ARLEN[1]       )
  ,.AXI_01_ARSIZE                (AXI_ARSIZE[1]      )
  ,.AXI_01_ARVALID               (AXI_ARVALID[1]     )
  ,.AXI_01_AWADDR                (AXI_AWADDR[1]      )
  ,.AXI_01_AWBURST               (AXI_AWBURST[1]     )
  ,.AXI_01_AWID                  (AXI_AWID[1]        )
  ,.AXI_01_AWLEN                 (AXI_AWLEN[1]       )
  ,.AXI_01_AWSIZE                (AXI_AWSIZE[1]      )
  ,.AXI_01_AWVALID               (AXI_AWVALID[1]     )
  ,.AXI_01_RREADY                (AXI_RREADY[1]      )
  ,.AXI_01_BREADY                (AXI_BREADY[1]      )
  ,.AXI_01_WDATA                 (AXI_WDATA[1]       )
  ,.AXI_01_WLAST                 (AXI_WLAST[1]       )
  ,.AXI_01_WSTRB                 (AXI_WSTRB[1]       )
  ,.AXI_01_WDATA_PARITY          (AXI_WDATA_PARITY[1])
  ,.AXI_01_WVALID                (AXI_WVALID[1]      )
  ,.AXI_02_ACLK                  (AXI_ACLK           )
  ,.AXI_02_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_02_ARADDR                (AXI_ARADDR[2]      )
  ,.AXI_02_ARBURST               (AXI_ARBURST[2]     )
  ,.AXI_02_ARID                  (AXI_ARID[2]        )
  ,.AXI_02_ARLEN                 (AXI_ARLEN[2]       )
  ,.AXI_02_ARSIZE                (AXI_ARSIZE[2]      )
  ,.AXI_02_ARVALID               (AXI_ARVALID[2]     )
  ,.AXI_02_AWADDR                (AXI_AWADDR[2]      )
  ,.AXI_02_AWBURST               (AXI_AWBURST[2]     )
  ,.AXI_02_AWID                  (AXI_AWID[2]        )
  ,.AXI_02_AWLEN                 (AXI_AWLEN[2]       )
  ,.AXI_02_AWSIZE                (AXI_AWSIZE[2]      )
  ,.AXI_02_AWVALID               (AXI_AWVALID[2]     )
  ,.AXI_02_RREADY                (AXI_RREADY[2]      )
  ,.AXI_02_BREADY                (AXI_BREADY[2]      )
  ,.AXI_02_WDATA                 (AXI_WDATA[2]       )
  ,.AXI_02_WLAST                 (AXI_WLAST[2]       )
  ,.AXI_02_WSTRB                 (AXI_WSTRB[2]       )
  ,.AXI_02_WDATA_PARITY          (AXI_WDATA_PARITY[2])
  ,.AXI_02_WVALID                (AXI_WVALID[2]      )
  ,.AXI_03_ACLK                  (AXI_ACLK           )
  ,.AXI_03_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_03_ARADDR                (AXI_ARADDR[3]      )
  ,.AXI_03_ARBURST               (AXI_ARBURST[3]     )
  ,.AXI_03_ARID                  (AXI_ARID[3]        )
  ,.AXI_03_ARLEN                 (AXI_ARLEN[3]       )
  ,.AXI_03_ARSIZE                (AXI_ARSIZE[3]      )
  ,.AXI_03_ARVALID               (AXI_ARVALID[3]     )
  ,.AXI_03_AWADDR                (AXI_AWADDR[3]      )
  ,.AXI_03_AWBURST               (AXI_AWBURST[3]     )
  ,.AXI_03_AWID                  (AXI_AWID[3]        )
  ,.AXI_03_AWLEN                 (AXI_AWLEN[3]       )
  ,.AXI_03_AWSIZE                (AXI_AWSIZE[3]      )
  ,.AXI_03_AWVALID               (AXI_AWVALID[3]     )
  ,.AXI_03_RREADY                (AXI_RREADY[3]      )
  ,.AXI_03_BREADY                (AXI_BREADY[3]      )
  ,.AXI_03_WDATA                 (AXI_WDATA[3]       )
  ,.AXI_03_WLAST                 (AXI_WLAST[3]       )
  ,.AXI_03_WSTRB                 (AXI_WSTRB[3]       )
  ,.AXI_03_WDATA_PARITY          (AXI_WDATA_PARITY[3])
  ,.AXI_03_WVALID                (AXI_WVALID[3]      )
  ,.AXI_04_ACLK                  (AXI_ACLK           )
  ,.AXI_04_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_04_ARADDR                (AXI_ARADDR[4]      )
  ,.AXI_04_ARBURST               (AXI_ARBURST[4]     )
  ,.AXI_04_ARID                  (AXI_ARID[4]        )
  ,.AXI_04_ARLEN                 (AXI_ARLEN[4]       )
  ,.AXI_04_ARSIZE                (AXI_ARSIZE[4]      )
  ,.AXI_04_ARVALID               (AXI_ARVALID[4]     )
  ,.AXI_04_AWADDR                (AXI_AWADDR[4]      )
  ,.AXI_04_AWBURST               (AXI_AWBURST[4]     )
  ,.AXI_04_AWID                  (AXI_AWID[4]        )
  ,.AXI_04_AWLEN                 (AXI_AWLEN[4]       )
  ,.AXI_04_AWSIZE                (AXI_AWSIZE[4]      )
  ,.AXI_04_AWVALID               (AXI_AWVALID[4]     )
  ,.AXI_04_RREADY                (AXI_RREADY[4]      )
  ,.AXI_04_BREADY                (AXI_BREADY[4]      )
  ,.AXI_04_WDATA                 (AXI_WDATA[4]       )
  ,.AXI_04_WLAST                 (AXI_WLAST[4]       )
  ,.AXI_04_WSTRB                 (AXI_WSTRB[4]       )
  ,.AXI_04_WDATA_PARITY          (AXI_WDATA_PARITY[4])
  ,.AXI_04_WVALID                (AXI_WVALID[4]      )
  ,.AXI_05_ACLK                  (AXI_ACLK           )
  ,.AXI_05_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_05_ARADDR                (AXI_ARADDR[5]      )
  ,.AXI_05_ARBURST               (AXI_ARBURST[5]     )
  ,.AXI_05_ARID                  (AXI_ARID[5]        )
  ,.AXI_05_ARLEN                 (AXI_ARLEN[5]       )
  ,.AXI_05_ARSIZE                (AXI_ARSIZE[5]      )
  ,.AXI_05_ARVALID               (AXI_ARVALID[5]     )
  ,.AXI_05_AWADDR                (AXI_AWADDR[5]      )
  ,.AXI_05_AWBURST               (AXI_AWBURST[5]     )
  ,.AXI_05_AWID                  (AXI_AWID[5]        )
  ,.AXI_05_AWLEN                 (AXI_AWLEN[5]       )
  ,.AXI_05_AWSIZE                (AXI_AWSIZE[5]      )
  ,.AXI_05_AWVALID               (AXI_AWVALID[5]     )
  ,.AXI_05_RREADY                (AXI_RREADY[5]      )
  ,.AXI_05_BREADY                (AXI_BREADY[5]      )
  ,.AXI_05_WDATA                 (AXI_WDATA[5]       )
  ,.AXI_05_WLAST                 (AXI_WLAST[5]       )
  ,.AXI_05_WSTRB                 (AXI_WSTRB[5]       )
  ,.AXI_05_WDATA_PARITY          (AXI_WDATA_PARITY[5])
  ,.AXI_05_WVALID                (AXI_WVALID[5]      )
  ,.AXI_06_ACLK                  (AXI_ACLK           )
  ,.AXI_06_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_06_ARADDR                (AXI_ARADDR[6]      )
  ,.AXI_06_ARBURST               (AXI_ARBURST[6]     )
  ,.AXI_06_ARID                  (AXI_ARID[6]        )
  ,.AXI_06_ARLEN                 (AXI_ARLEN[6]       )
  ,.AXI_06_ARSIZE                (AXI_ARSIZE[6]      )
  ,.AXI_06_ARVALID               (AXI_ARVALID[6]     )
  ,.AXI_06_AWADDR                (AXI_AWADDR[6]      )
  ,.AXI_06_AWBURST               (AXI_AWBURST[6]     )
  ,.AXI_06_AWID                  (AXI_AWID[6]        )
  ,.AXI_06_AWLEN                 (AXI_AWLEN[6]       )
  ,.AXI_06_AWSIZE                (AXI_AWSIZE[6]      )
  ,.AXI_06_AWVALID               (AXI_AWVALID[6]     )
  ,.AXI_06_RREADY                (AXI_RREADY[6]      )
  ,.AXI_06_BREADY                (AXI_BREADY[6]      )
  ,.AXI_06_WDATA                 (AXI_WDATA[6]       )
  ,.AXI_06_WLAST                 (AXI_WLAST[6]       )
  ,.AXI_06_WSTRB                 (AXI_WSTRB[6]       )
  ,.AXI_06_WDATA_PARITY          (AXI_WDATA_PARITY[6])
  ,.AXI_06_WVALID                (AXI_WVALID[6]      )
  ,.AXI_07_ACLK                  (AXI_ACLK           )
  ,.AXI_07_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_07_ARADDR                (AXI_ARADDR[7]      )
  ,.AXI_07_ARBURST               (AXI_ARBURST[7]     )
  ,.AXI_07_ARID                  (AXI_ARID[7]        )
  ,.AXI_07_ARLEN                 (AXI_ARLEN[7]       )
  ,.AXI_07_ARSIZE                (AXI_ARSIZE[7]      )
  ,.AXI_07_ARVALID               (AXI_ARVALID[7]     )
  ,.AXI_07_AWADDR                (AXI_AWADDR[7]      )
  ,.AXI_07_AWBURST               (AXI_AWBURST[7]     )
  ,.AXI_07_AWID                  (AXI_AWID[7]        )
  ,.AXI_07_AWLEN                 (AXI_AWLEN[7]       )
  ,.AXI_07_AWSIZE                (AXI_AWSIZE[7]      )
  ,.AXI_07_AWVALID               (AXI_AWVALID[7]     )
  ,.AXI_07_RREADY                (AXI_RREADY[7]      )
  ,.AXI_07_BREADY                (AXI_BREADY[7]      )
  ,.AXI_07_WDATA                 (AXI_WDATA[7]       )
  ,.AXI_07_WLAST                 (AXI_WLAST[7]       )
  ,.AXI_07_WSTRB                 (AXI_WSTRB[7]       )
  ,.AXI_07_WDATA_PARITY          (AXI_WDATA_PARITY[7])
  ,.AXI_07_WVALID                (AXI_WVALID[7]      )
  ,.AXI_08_ACLK                  (AXI_ACLK           )
  ,.AXI_08_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_08_ARADDR                (AXI_ARADDR[8]      )
  ,.AXI_08_ARBURST               (AXI_ARBURST[8]     )
  ,.AXI_08_ARID                  (AXI_ARID[8]        )
  ,.AXI_08_ARLEN                 (AXI_ARLEN[8]       )
  ,.AXI_08_ARSIZE                (AXI_ARSIZE[8]      )
  ,.AXI_08_ARVALID               (AXI_ARVALID[8]     )
  ,.AXI_08_AWADDR                (AXI_AWADDR[8]      )
  ,.AXI_08_AWBURST               (AXI_AWBURST[8]     )
  ,.AXI_08_AWID                  (AXI_AWID[8]        )
  ,.AXI_08_AWLEN                 (AXI_AWLEN[8]       )
  ,.AXI_08_AWSIZE                (AXI_AWSIZE[8]      )
  ,.AXI_08_AWVALID               (AXI_AWVALID[8]     )
  ,.AXI_08_RREADY                (AXI_RREADY[8]      )
  ,.AXI_08_BREADY                (AXI_BREADY[8]      )
  ,.AXI_08_WDATA                 (AXI_WDATA[8]       )
  ,.AXI_08_WLAST                 (AXI_WLAST[8]       )
  ,.AXI_08_WSTRB                 (AXI_WSTRB[8]       )
  ,.AXI_08_WDATA_PARITY          (AXI_WDATA_PARITY[8])
  ,.AXI_08_WVALID                (AXI_WVALID[8]      )
  ,.AXI_09_ACLK                  (AXI_ACLK           )
  ,.AXI_09_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_09_ARADDR                (AXI_ARADDR[9]      )
  ,.AXI_09_ARBURST               (AXI_ARBURST[9]     )
  ,.AXI_09_ARID                  (AXI_ARID[9]        )
  ,.AXI_09_ARLEN                 (AXI_ARLEN[9]       )
  ,.AXI_09_ARSIZE                (AXI_ARSIZE[9]      )
  ,.AXI_09_ARVALID               (AXI_ARVALID[9]     )
  ,.AXI_09_AWADDR                (AXI_AWADDR[9]      )
  ,.AXI_09_AWBURST               (AXI_AWBURST[9]     )
  ,.AXI_09_AWID                  (AXI_AWID[9]        )
  ,.AXI_09_AWLEN                 (AXI_AWLEN[9]       )
  ,.AXI_09_AWSIZE                (AXI_AWSIZE[9]      )
  ,.AXI_09_AWVALID               (AXI_AWVALID[9]     )
  ,.AXI_09_RREADY                (AXI_RREADY[9]      )
  ,.AXI_09_BREADY                (AXI_BREADY[9]      )
  ,.AXI_09_WDATA                 (AXI_WDATA[9]       )
  ,.AXI_09_WLAST                 (AXI_WLAST[9]       )
  ,.AXI_09_WSTRB                 (AXI_WSTRB[9]       )
  ,.AXI_09_WDATA_PARITY          (AXI_WDATA_PARITY[9])
  ,.AXI_09_WVALID                (AXI_WVALID[9]      )
  ,.AXI_10_ACLK                  (AXI_ACLK           )
  ,.AXI_10_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_10_ARADDR                (AXI_ARADDR[10]      )
  ,.AXI_10_ARBURST               (AXI_ARBURST[10]     )
  ,.AXI_10_ARID                  (AXI_ARID[10]        )
  ,.AXI_10_ARLEN                 (AXI_ARLEN[10]       )
  ,.AXI_10_ARSIZE                (AXI_ARSIZE[10]      )
  ,.AXI_10_ARVALID               (AXI_ARVALID[10]     )
  ,.AXI_10_AWADDR                (AXI_AWADDR[10]      )
  ,.AXI_10_AWBURST               (AXI_AWBURST[10]     )
  ,.AXI_10_AWID                  (AXI_AWID[10]        )
  ,.AXI_10_AWLEN                 (AXI_AWLEN[10]       )
  ,.AXI_10_AWSIZE                (AXI_AWSIZE[10]      )
  ,.AXI_10_AWVALID               (AXI_AWVALID[10]     )
  ,.AXI_10_RREADY                (AXI_RREADY[10]      )
  ,.AXI_10_BREADY                (AXI_BREADY[10]      )
  ,.AXI_10_WDATA                 (AXI_WDATA[10]       )
  ,.AXI_10_WLAST                 (AXI_WLAST[10]       )
  ,.AXI_10_WSTRB                 (AXI_WSTRB[10]       )
  ,.AXI_10_WDATA_PARITY          (AXI_WDATA_PARITY[10])
  ,.AXI_10_WVALID                (AXI_WVALID[10]      )
  ,.AXI_11_ACLK                  (AXI_ACLK           )
  ,.AXI_11_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_11_ARADDR                (AXI_ARADDR[11]      )
  ,.AXI_11_ARBURST               (AXI_ARBURST[11]     )
  ,.AXI_11_ARID                  (AXI_ARID[11]        )
  ,.AXI_11_ARLEN                 (AXI_ARLEN[11]       )
  ,.AXI_11_ARSIZE                (AXI_ARSIZE[11]      )
  ,.AXI_11_ARVALID               (AXI_ARVALID[11]     )
  ,.AXI_11_AWADDR                (AXI_AWADDR[11]      )
  ,.AXI_11_AWBURST               (AXI_AWBURST[11]     )
  ,.AXI_11_AWID                  (AXI_AWID[11]        )
  ,.AXI_11_AWLEN                 (AXI_AWLEN[11]       )
  ,.AXI_11_AWSIZE                (AXI_AWSIZE[11]      )
  ,.AXI_11_AWVALID               (AXI_AWVALID[11]     )
  ,.AXI_11_RREADY                (AXI_RREADY[11]      )
  ,.AXI_11_BREADY                (AXI_BREADY[11]      )
  ,.AXI_11_WDATA                 (AXI_WDATA[11]       )
  ,.AXI_11_WLAST                 (AXI_WLAST[11]       )
  ,.AXI_11_WSTRB                 (AXI_WSTRB[11]       )
  ,.AXI_11_WDATA_PARITY          (AXI_WDATA_PARITY[11])
  ,.AXI_11_WVALID                (AXI_WVALID[11]      )
  ,.AXI_12_ACLK                  (AXI_ACLK           )
  ,.AXI_12_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_12_ARADDR                (AXI_ARADDR[12]      )
  ,.AXI_12_ARBURST               (AXI_ARBURST[12]     )
  ,.AXI_12_ARID                  (AXI_ARID[12]        )
  ,.AXI_12_ARLEN                 (AXI_ARLEN[12]       )
  ,.AXI_12_ARSIZE                (AXI_ARSIZE[12]      )
  ,.AXI_12_ARVALID               (AXI_ARVALID[12]     )
  ,.AXI_12_AWADDR                (AXI_AWADDR[12]      )
  ,.AXI_12_AWBURST               (AXI_AWBURST[12]     )
  ,.AXI_12_AWID                  (AXI_AWID[12]        )
  ,.AXI_12_AWLEN                 (AXI_AWLEN[12]       )
  ,.AXI_12_AWSIZE                (AXI_AWSIZE[12]      )
  ,.AXI_12_AWVALID               (AXI_AWVALID[12]     )
  ,.AXI_12_RREADY                (AXI_RREADY[12]      )
  ,.AXI_12_BREADY                (AXI_BREADY[12]      )
  ,.AXI_12_WDATA                 (AXI_WDATA[12]       )
  ,.AXI_12_WLAST                 (AXI_WLAST[12]       )
  ,.AXI_12_WSTRB                 (AXI_WSTRB[12]       )
  ,.AXI_12_WDATA_PARITY          (AXI_WDATA_PARITY[12])
  ,.AXI_12_WVALID                (AXI_WVALID[12]      )
  ,.AXI_13_ACLK                  (AXI_ACLK           )
  ,.AXI_13_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_13_ARADDR                (AXI_ARADDR[13]      )
  ,.AXI_13_ARBURST               (AXI_ARBURST[13]     )
  ,.AXI_13_ARID                  (AXI_ARID[13]        )
  ,.AXI_13_ARLEN                 (AXI_ARLEN[13]       )
  ,.AXI_13_ARSIZE                (AXI_ARSIZE[13]      )
  ,.AXI_13_ARVALID               (AXI_ARVALID[13]     )
  ,.AXI_13_AWADDR                (AXI_AWADDR[13]      )
  ,.AXI_13_AWBURST               (AXI_AWBURST[13]     )
  ,.AXI_13_AWID                  (AXI_AWID[13]        )
  ,.AXI_13_AWLEN                 (AXI_AWLEN[13]       )
  ,.AXI_13_AWSIZE                (AXI_AWSIZE[13]      )
  ,.AXI_13_AWVALID               (AXI_AWVALID[13]     )
  ,.AXI_13_RREADY                (AXI_RREADY[13]      )
  ,.AXI_13_BREADY                (AXI_BREADY[13]      )
  ,.AXI_13_WDATA                 (AXI_WDATA[13]       )
  ,.AXI_13_WLAST                 (AXI_WLAST[13]       )
  ,.AXI_13_WSTRB                 (AXI_WSTRB[13]       )
  ,.AXI_13_WDATA_PARITY          (AXI_WDATA_PARITY[13])
  ,.AXI_13_WVALID                (AXI_WVALID[13]      )
  ,.AXI_14_ACLK                  (AXI_ACLK           )
  ,.AXI_14_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_14_ARADDR                (AXI_ARADDR[14]      )
  ,.AXI_14_ARBURST               (AXI_ARBURST[14]     )
  ,.AXI_14_ARID                  (AXI_ARID[14]        )
  ,.AXI_14_ARLEN                 (AXI_ARLEN[14]       )
  ,.AXI_14_ARSIZE                (AXI_ARSIZE[14]      )
  ,.AXI_14_ARVALID               (AXI_ARVALID[14]     )
  ,.AXI_14_AWADDR                (AXI_AWADDR[14]      )
  ,.AXI_14_AWBURST               (AXI_AWBURST[14]     )
  ,.AXI_14_AWID                  (AXI_AWID[14]        )
  ,.AXI_14_AWLEN                 (AXI_AWLEN[14]       )
  ,.AXI_14_AWSIZE                (AXI_AWSIZE[14]      )
  ,.AXI_14_AWVALID               (AXI_AWVALID[14]     )
  ,.AXI_14_RREADY                (AXI_RREADY[14]      )
  ,.AXI_14_BREADY                (AXI_BREADY[14]      )
  ,.AXI_14_WDATA                 (AXI_WDATA[14]       )
  ,.AXI_14_WLAST                 (AXI_WLAST[14]       )
  ,.AXI_14_WSTRB                 (AXI_WSTRB[14]       )
  ,.AXI_14_WDATA_PARITY          (AXI_WDATA_PARITY[14])
  ,.AXI_14_WVALID                (AXI_WVALID[14]      )
  ,.AXI_15_ACLK                  (AXI_ACLK           )
  ,.AXI_15_ARESET_N              (AXI_ARESET_N       )
  ,.AXI_15_ARADDR                (AXI_ARADDR[15]      )
  ,.AXI_15_ARBURST               (AXI_ARBURST[15]     )
  ,.AXI_15_ARID                  (AXI_ARID[15]        )
  ,.AXI_15_ARLEN                 (AXI_ARLEN[15]       )
  ,.AXI_15_ARSIZE                (AXI_ARSIZE[15]      )
  ,.AXI_15_ARVALID               (AXI_ARVALID[15]     )
  ,.AXI_15_AWADDR                (AXI_AWADDR[15]      )
  ,.AXI_15_AWBURST               (AXI_AWBURST[15]     )
  ,.AXI_15_AWID                  (AXI_AWID[15]        )
  ,.AXI_15_AWLEN                 (AXI_AWLEN[15]       )
  ,.AXI_15_AWSIZE                (AXI_AWSIZE[15]      )
  ,.AXI_15_AWVALID               (AXI_AWVALID[15]     )
  ,.AXI_15_RREADY                (AXI_RREADY[15]      )
  ,.AXI_15_BREADY                (AXI_BREADY[15]      )
  ,.AXI_15_WDATA                 (AXI_WDATA[15]       )
  ,.AXI_15_WLAST                 (AXI_WLAST[15]       )
  ,.AXI_15_WSTRB                 (AXI_WSTRB[15]       )
  ,.AXI_15_WDATA_PARITY          (AXI_WDATA_PARITY[15])
  ,.AXI_15_WVALID                (AXI_WVALID[15]      )

  ,.APB_0_PCLK                   (APB_0_PCLK    )
  ,.APB_0_PRESET_N               (APB_hbm_reset)
  ,.APB_0_PWDATA                 (APB_0_PWDATA  )
  ,.APB_0_PADDR                  (APB_0_PADDR   )
  ,.APB_0_PENABLE                (APB_0_PENABLE )
  ,.APB_0_PSEL                   (APB_0_PSEL    )
  ,.APB_0_PWRITE                 (APB_0_PWRITE  )
  
  ,.AXI_00_ARREADY               (AXI_ARREADY[0]     )
  ,.AXI_00_AWREADY               (AXI_AWREADY[0]     )
  ,.AXI_00_RDATA_PARITY          (AXI_RDATA_PARITY[0])
  ,.AXI_00_RDATA                 (AXI_RDATA[0]       )
  ,.AXI_00_RID                   (AXI_RID[0]         )
  ,.AXI_00_RLAST                 (AXI_RLAST[0]       )
  ,.AXI_00_RRESP                 (AXI_RRESP[0]       )
  ,.AXI_00_RVALID                (AXI_RVALID[0]      )
  ,.AXI_00_WREADY                (AXI_WREADY[0]      )
  ,.AXI_00_BID                   (AXI_BID[0]         )
  ,.AXI_00_BRESP                 (AXI_BRESP[0]       )
  ,.AXI_00_BVALID                (AXI_BVALID[0]      )
  ,.AXI_01_ARREADY               (AXI_ARREADY[1]     )
  ,.AXI_01_AWREADY               (AXI_AWREADY[1]     )
  ,.AXI_01_RDATA_PARITY          (AXI_RDATA_PARITY[1])
  ,.AXI_01_RDATA                 (AXI_RDATA[1]       )
  ,.AXI_01_RID                   (AXI_RID[1]         )
  ,.AXI_01_RLAST                 (AXI_RLAST[1]       )
  ,.AXI_01_RRESP                 (AXI_RRESP[1]       )
  ,.AXI_01_RVALID                (AXI_RVALID[1]      )
  ,.AXI_01_WREADY                (AXI_WREADY[1]      )
  ,.AXI_01_BID                   (AXI_BID[1]         )
  ,.AXI_01_BRESP                 (AXI_BRESP[1]       )
  ,.AXI_01_BVALID                (AXI_BVALID[1]      )
  ,.AXI_02_ARREADY               (AXI_ARREADY[2]     )
  ,.AXI_02_AWREADY               (AXI_AWREADY[2]     )
  ,.AXI_02_RDATA_PARITY          (AXI_RDATA_PARITY[2])
  ,.AXI_02_RDATA                 (AXI_RDATA[2]       )
  ,.AXI_02_RID                   (AXI_RID[2]         )
  ,.AXI_02_RLAST                 (AXI_RLAST[2]       )
  ,.AXI_02_RRESP                 (AXI_RRESP[2]       )
  ,.AXI_02_RVALID                (AXI_RVALID[2]      )
  ,.AXI_02_WREADY                (AXI_WREADY[2]      )
  ,.AXI_02_BID                   (AXI_BID[2]         )
  ,.AXI_02_BRESP                 (AXI_BRESP[2]       )
  ,.AXI_02_BVALID                (AXI_BVALID[2]      )
  ,.AXI_03_ARREADY               (AXI_ARREADY[3]     )
  ,.AXI_03_AWREADY               (AXI_AWREADY[3]     )
  ,.AXI_03_RDATA_PARITY          (AXI_RDATA_PARITY[3])
  ,.AXI_03_RDATA                 (AXI_RDATA[3]       )
  ,.AXI_03_RID                   (AXI_RID[3]         )
  ,.AXI_03_RLAST                 (AXI_RLAST[3]       )
  ,.AXI_03_RRESP                 (AXI_RRESP[3]       )
  ,.AXI_03_RVALID                (AXI_RVALID[3]      )
  ,.AXI_03_WREADY                (AXI_WREADY[3]      )
  ,.AXI_03_BID                   (AXI_BID[3]         )
  ,.AXI_03_BRESP                 (AXI_BRESP[3]       )
  ,.AXI_03_BVALID                (AXI_BVALID[3]      )
  ,.AXI_04_ARREADY               (AXI_ARREADY[4]     )
  ,.AXI_04_AWREADY               (AXI_AWREADY[4]     )
  ,.AXI_04_RDATA_PARITY          (AXI_RDATA_PARITY[4])
  ,.AXI_04_RDATA                 (AXI_RDATA[4]       )
  ,.AXI_04_RID                   (AXI_RID[4]         )
  ,.AXI_04_RLAST                 (AXI_RLAST[4]       )
  ,.AXI_04_RRESP                 (AXI_RRESP[4]       )
  ,.AXI_04_RVALID                (AXI_RVALID[4]      )
  ,.AXI_04_WREADY                (AXI_WREADY[4]      )
  ,.AXI_04_BID                   (AXI_BID[4]         )
  ,.AXI_04_BRESP                 (AXI_BRESP[4]       )
  ,.AXI_04_BVALID                (AXI_BVALID[4]      )
  ,.AXI_05_ARREADY               (AXI_ARREADY[5]     )
  ,.AXI_05_AWREADY               (AXI_AWREADY[5]     )
  ,.AXI_05_RDATA_PARITY          (AXI_RDATA_PARITY[5])
  ,.AXI_05_RDATA                 (AXI_RDATA[5]       )
  ,.AXI_05_RID                   (AXI_RID[5]         )
  ,.AXI_05_RLAST                 (AXI_RLAST[5]       )
  ,.AXI_05_RRESP                 (AXI_RRESP[5]       )
  ,.AXI_05_RVALID                (AXI_RVALID[5]      )
  ,.AXI_05_WREADY                (AXI_WREADY[5]      )
  ,.AXI_05_BID                   (AXI_BID[5]         )
  ,.AXI_05_BRESP                 (AXI_BRESP[5]       )
  ,.AXI_05_BVALID                (AXI_BVALID[5]      )
  ,.AXI_06_ARREADY               (AXI_ARREADY[6]     )
  ,.AXI_06_AWREADY               (AXI_AWREADY[6]     )
  ,.AXI_06_RDATA_PARITY          (AXI_RDATA_PARITY[6])
  ,.AXI_06_RDATA                 (AXI_RDATA[6]       )
  ,.AXI_06_RID                   (AXI_RID[6]         )
  ,.AXI_06_RLAST                 (AXI_RLAST[6]       )
  ,.AXI_06_RRESP                 (AXI_RRESP[6]       )
  ,.AXI_06_RVALID                (AXI_RVALID[6]      )
  ,.AXI_06_WREADY                (AXI_WREADY[6]      )
  ,.AXI_06_BID                   (AXI_BID[6]         )
  ,.AXI_06_BRESP                 (AXI_BRESP[6]       )
  ,.AXI_06_BVALID                (AXI_BVALID[6]      )
  ,.AXI_07_ARREADY               (AXI_ARREADY[7]     )
  ,.AXI_07_AWREADY               (AXI_AWREADY[7]     )
  ,.AXI_07_RDATA_PARITY          (AXI_RDATA_PARITY[7])
  ,.AXI_07_RDATA                 (AXI_RDATA[7]       )
  ,.AXI_07_RID                   (AXI_RID[7]         )
  ,.AXI_07_RLAST                 (AXI_RLAST[7]       )
  ,.AXI_07_RRESP                 (AXI_RRESP[7]       )
  ,.AXI_07_RVALID                (AXI_RVALID[7]      )
  ,.AXI_07_WREADY                (AXI_WREADY[7]      )
  ,.AXI_07_BID                   (AXI_BID[7]         )
  ,.AXI_07_BRESP                 (AXI_BRESP[7]       )
  ,.AXI_07_BVALID                (AXI_BVALID[7]      )
  ,.AXI_08_ARREADY               (AXI_ARREADY[8]     )
  ,.AXI_08_AWREADY               (AXI_AWREADY[8]     )
  ,.AXI_08_RDATA_PARITY          (AXI_RDATA_PARITY[8])
  ,.AXI_08_RDATA                 (AXI_RDATA[8]       )
  ,.AXI_08_RID                   (AXI_RID[8]         )
  ,.AXI_08_RLAST                 (AXI_RLAST[8]       )
  ,.AXI_08_RRESP                 (AXI_RRESP[8]       )
  ,.AXI_08_RVALID                (AXI_RVALID[8]      )
  ,.AXI_08_WREADY                (AXI_WREADY[8]      )
  ,.AXI_08_BID                   (AXI_BID[8]         )
  ,.AXI_08_BRESP                 (AXI_BRESP[8]       )
  ,.AXI_08_BVALID                (AXI_BVALID[8]      )
  ,.AXI_09_ARREADY               (AXI_ARREADY[9]     )
  ,.AXI_09_AWREADY               (AXI_AWREADY[9]     )
  ,.AXI_09_RDATA_PARITY          (AXI_RDATA_PARITY[9])
  ,.AXI_09_RDATA                 (AXI_RDATA[9]       )
  ,.AXI_09_RID                   (AXI_RID[9]         )
  ,.AXI_09_RLAST                 (AXI_RLAST[9]       )
  ,.AXI_09_RRESP                 (AXI_RRESP[9]       )
  ,.AXI_09_RVALID                (AXI_RVALID[9]      )
  ,.AXI_09_WREADY                (AXI_WREADY[9]      )
  ,.AXI_09_BID                   (AXI_BID[9]         )
  ,.AXI_09_BRESP                 (AXI_BRESP[9]       )
  ,.AXI_09_BVALID                (AXI_BVALID[9]      )
  ,.AXI_10_ARREADY               (AXI_ARREADY[10]     )
  ,.AXI_10_AWREADY               (AXI_AWREADY[10]     )
  ,.AXI_10_RDATA_PARITY          (AXI_RDATA_PARITY[10])
  ,.AXI_10_RDATA                 (AXI_RDATA[10]       )
  ,.AXI_10_RID                   (AXI_RID[10]         )
  ,.AXI_10_RLAST                 (AXI_RLAST[10]       )
  ,.AXI_10_RRESP                 (AXI_RRESP[10]       )
  ,.AXI_10_RVALID                (AXI_RVALID[10]      )
  ,.AXI_10_WREADY                (AXI_WREADY[10]      )
  ,.AXI_10_BID                   (AXI_BID[10]         )
  ,.AXI_10_BRESP                 (AXI_BRESP[10]       )
  ,.AXI_10_BVALID                (AXI_BVALID[10]      )
  ,.AXI_11_ARREADY               (AXI_ARREADY[11]     )
  ,.AXI_11_AWREADY               (AXI_AWREADY[11]     )
  ,.AXI_11_RDATA_PARITY          (AXI_RDATA_PARITY[11])
  ,.AXI_11_RDATA                 (AXI_RDATA[11]       )
  ,.AXI_11_RID                   (AXI_RID[11]         )
  ,.AXI_11_RLAST                 (AXI_RLAST[11]       )
  ,.AXI_11_RRESP                 (AXI_RRESP[11]       )
  ,.AXI_11_RVALID                (AXI_RVALID[11]      )
  ,.AXI_11_WREADY                (AXI_WREADY[11]      )
  ,.AXI_11_BID                   (AXI_BID[11]         )
  ,.AXI_11_BRESP                 (AXI_BRESP[11]       )
  ,.AXI_11_BVALID                (AXI_BVALID[11]      )
  ,.AXI_12_ARREADY               (AXI_ARREADY[12]     )
  ,.AXI_12_AWREADY               (AXI_AWREADY[12]     )
  ,.AXI_12_RDATA_PARITY          (AXI_RDATA_PARITY[12])
  ,.AXI_12_RDATA                 (AXI_RDATA[12]       )
  ,.AXI_12_RID                   (AXI_RID[12]         )
  ,.AXI_12_RLAST                 (AXI_RLAST[12]       )
  ,.AXI_12_RRESP                 (AXI_RRESP[12]       )
  ,.AXI_12_RVALID                (AXI_RVALID[12]      )
  ,.AXI_12_WREADY                (AXI_WREADY[12]      )
  ,.AXI_12_BID                   (AXI_BID[12]         )
  ,.AXI_12_BRESP                 (AXI_BRESP[12]       )
  ,.AXI_12_BVALID                (AXI_BVALID[12]      )
  ,.AXI_13_ARREADY               (AXI_ARREADY[13]     )
  ,.AXI_13_AWREADY               (AXI_AWREADY[13]     )
  ,.AXI_13_RDATA_PARITY          (AXI_RDATA_PARITY[13])
  ,.AXI_13_RDATA                 (AXI_RDATA[13]       )
  ,.AXI_13_RID                   (AXI_RID[13]         )
  ,.AXI_13_RLAST                 (AXI_RLAST[13]       )
  ,.AXI_13_RRESP                 (AXI_RRESP[13]       )
  ,.AXI_13_RVALID                (AXI_RVALID[13]      )
  ,.AXI_13_WREADY                (AXI_WREADY[13]      )
  ,.AXI_13_BID                   (AXI_BID[13]         )
  ,.AXI_13_BRESP                 (AXI_BRESP[13]       )
  ,.AXI_13_BVALID                (AXI_BVALID[13]      )
  ,.AXI_14_ARREADY               (AXI_ARREADY[14]     )
  ,.AXI_14_AWREADY               (AXI_AWREADY[14]     )
  ,.AXI_14_RDATA_PARITY          (AXI_RDATA_PARITY[14])
  ,.AXI_14_RDATA                 (AXI_RDATA[14]       )
  ,.AXI_14_RID                   (AXI_RID[14]         )
  ,.AXI_14_RLAST                 (AXI_RLAST[14]       )
  ,.AXI_14_RRESP                 (AXI_RRESP[14]       )
  ,.AXI_14_RVALID                (AXI_RVALID[14]      )
  ,.AXI_14_WREADY                (AXI_WREADY[14]      )
  ,.AXI_14_BID                   (AXI_BID[14]         )
  ,.AXI_14_BRESP                 (AXI_BRESP[14]       )
  ,.AXI_14_BVALID                (AXI_BVALID[14]      )
  ,.AXI_15_ARREADY               (AXI_ARREADY[15]     )
  ,.AXI_15_AWREADY               (AXI_AWREADY[15]     )
  ,.AXI_15_RDATA_PARITY          (AXI_RDATA_PARITY[15])
  ,.AXI_15_RDATA                 (AXI_RDATA[15]       )
  ,.AXI_15_RID                   (AXI_RID[15]         )
  ,.AXI_15_RLAST                 (AXI_RLAST[15]       )
  ,.AXI_15_RRESP                 (AXI_RRESP[15]       )
  ,.AXI_15_RVALID                (AXI_RVALID[15]      )
  ,.AXI_15_WREADY                (AXI_WREADY[15]      )
  ,.AXI_15_BID                   (AXI_BID[15]         )
  ,.AXI_15_BRESP                 (AXI_BRESP[15]       )
  ,.AXI_15_BVALID                (AXI_BVALID[15]      )
  ,.apb_complete_0               (apb_complete_0)
  ,.APB_0_PRDATA                 (APB_0_PRDATA )
  ,.APB_0_PREADY                 (APB_0_PREADY )
  ,.APB_0_PSLVERR                (APB_0_PSLVERR)
  
  ,.DRAM_0_STAT_CATTRIP          ()
  ,.DRAM_0_STAT_TEMP             ()
);
	
endmodule
